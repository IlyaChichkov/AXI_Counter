module m_axi_reg
(

);

logic crc_module_en;

endmodule